module wave_display (
    input clk,
    input reset,
    input [10:0] x,  // [0..1279]
    input [9:0]  y,  // [0..1023]
    input valid,
    input [7:0] read_value,
    input read_index,
    output wire [8:0] read_address,
    output wire valid_pixel,
    output wire [7:0] r,
    output wire [7:0] g,
    output wire [7:0] b
);

//read address: concat read index, x[9], then 7 bits of x not counting lsb
assign read_address = {read_index, x[9], x[7:1]};
	
//adjust for aspect ratio/screen size
wire [7:0] read_value_adjusted = (read_value >> 1) + 8'd32;

//take 8:1 bits of y for the y value
wire [7:0] y_val;
assign y_val = y[8:1];
//pixel is valid if 9th and 8th bit is 01 or 10, so we use xor. also, clip the top y-vals to get rid of artifacts
assign valid_pixel = ((x[10:9] == 2'b01) || (x[10:9] == 2'b0)) & valid & (x > 11'b00100000010);


//FFs
wire [8:0] prev_addr;
dffr #(9) read_addr_ff(
	.clk(clk), 
	.r(reset), 
	.d(read_address), 
	.q(prev_addr));
wire [7:0] prev_value;
dffre #(8) read_value_ff(
	.clk(clk), 
	.r(reset), 
	.en(read_address != prev_addr), 
	.d(read_value_adjusted), 
	.q(prev_value));

//when to display: between min and max of cur and prev y val
reg display;
always @(*) begin
	if(y_val >= prev_value && y_val <= read_value_adjusted) display = 1; //prev_value < read_value
	else if(y_val <= prev_value && y_val >= read_value_adjusted) display = 1; //prev_value > read_value
	else display = 0;
end

assign {r,g,b} = (display & valid) ? 24'hFFFFFF : 24'h000000;
endmodule
